module addr2b_hex8seg_EGo1(
)