module and21(D0,D1,Y);

	input D0;
	input D1;
	output Y;

	wire D0,D1,Y;

	assign Y = D0 & D1;

endmodule